/// # parsing
open sm'_operators

/// ## fparsec

/// ## parsing

/// ### position

/// ### range
type range =
    {
        from : int
        to : int
    }

type position =
    {
        line : int
        col : int
    }

/// ### parser_state
nominal parser_state =
    {
        line_text : sm'.string_builder
        position : position
    }

/// ### new_parser_state
inl new_parser_state line_text (line : i32) (col : i32) =
    { line_text = line_text |> sm'.string_builder; position = { line col } }

/// ### new_parser_state'
inl new_parser_state' () =
    new_parser_state "" 1 1 |> parser_state

/// ### parser
type parser t = string * int * parser_state -> result (t * int * parser_state) string

/// ### parse
inl parse forall t.
    (p : parser t)
    (input : string)
    (s : parser_state)
    : result (t * string * parser_state) string
    =
    p (input, 0, s)
    |> resultm.map fun result, i, s' =>
        result,
        input |> sm'.range (am'.Start i) (am'.End eval),
        s'

/// ### inc
inl inc (parser_state s) = function
    | '\n' => { line = s.position.line + 1; col = 1 }
    | _ => { s.position with col = s.position.col + 1 }.position

/// ### update_char
inl update_char (parser_state s as s') (c : char) : parser_state =
    { s with
        position =
            match c with
            | '\n' => { line = s.position.line + 1; col = 1 }
            | _ => { s.position with col = s.position.col + 1 }.position
        line_text =
            match c with
            | '\n' => s.line_text |> sm'.builder_clear
            | _ => s.line_text |> sm'.builder_append $c
    } |> parser_state

/// ### update
inl update result s =
    let rec 루프 (i : int) s =
        if i >= (result |> sm'.length)
        then s
        else result |> sm'.index i |> update_char s |> 루프 (i + 1)
    s |> 루프 0

/// ### run_parser
inl run_parser parser input =
    input
    |> parse parser
    |> fun parser => parser (new_parser_state' ())

/// ### any_char
inl any_char () : parser char = fun input, i, s =>
    if i >= (input |> sm'.length)
    then "parsing.any_char / unexpected end of input / " ++# ({ s } |> sm'.format) |> Error
    else
        inl c = input |> sm'.index i
        Ok (c, i + 1, c |> update_char s)

/// ### get_max_context
inl get_max_context () =
    120

/// ### p_char
inl p_char (c : char) : parser char =
    fun input, i, (parser_state ({ line_text position = { line col } } as s) as s') =>
        if i >= (input |> sm'.length)
        then "parsing.p_char / unexpected end of input / " ++# ({ c s } |> sm'.format) |> Error
        else
            inl got = input |> sm'.index i
            if got = c
            then Ok (got, i + 1, got |> update_char s')
            else
                inl total_len = input |> sm'.length
                inl end_line =
                    match input |> sm'.index_of_char_from i '\n' with
                    | -1 => total_len
                    | j  => (if j >= i then j else i + j) |> min total_len
                inl end = (i + get_max_context ()) |> min end_line |> min total_len
                inl rest = input |> sm'.range (am'.Start i) (am'.End fun _ => end)
                inl pointer_line = (" " |> sm'.replicate (col - 1)) ++# "^"
                "parsing.p_char / "
                ++# ({ expected = c; line col } |> sm'.format)
                ++# "\n" ++# $line_text ++# rest
                ++# "\n" ++# pointer_line ++# "\n"
                |> Error

/// ### any_string
inl any_string length : parser string = fun input, i, s =>
    if (input |> sm'.length) - i < length
    then "parsing.any_string / unexpected end of input / " ++# ({ s } |> sm'.format) |> Error
    else
        inl result = input |> sm'.range (am'.Start i) (am'.End fun _ => i + length)
        Ok (
            result,
            i + length,
            s |> update result
        )

/// ### skip_any_string
inl skip_any_string length : parser () = fun input, i, s =>
    if (input |> sm'.length) - i < length
    then "parsing.skip_any_string / unexpected end of input / " ++# ({ s } |> sm'.format) |> Error
    else
        Ok (
            (),
            i + length,
            s |> update (input |> sm'.range (am'.Start i) (am'.End fun _ => i + length))
        )

/// ### (>>.)
inl (>>.) forall t u. (a : parser t) (b : parser u) : parser u = fun input, i, s =>
    match a (input, i, s) with
    | Ok (_, i', s') => b (input, i', s')
    | Error e => Error e

/// ### (>>.)
inl (.>>) forall t u. (a : parser t) (b : parser u) : parser t = fun input, i, s =>
    match a (input, i, s) with
    | Ok (ra, i', s') =>
        b (input, i', s')
        |> resultm.map fun _, i'', s'' =>
            ra, i'', s''
    | Error e => Error e

/// ### (.>>.)
inl (.>>.) forall t u. (a : parser t) (b : parser u) : parser (t * u) = fun input, i, s =>
    match a (input, i, s) with
    | Ok (ra, i', s') =>
        b (input,  i', s')
        |> resultm.map fun rb, i'', s'' =>
            (ra, rb), i'', s''
    | Error e => Error e

/// ### (>>%)
inl (>>%) forall t u. (a : parser t) (b : u) : parser u =
    a >> resultm.map fun _, i', s' =>
        b, i', s'

/// ### none_of
inl none_of (chars : list char) : parser char = fun input, i, s =>
    inl chars' () : string =
        backend_switch {
            Gleam = fun () => chars |> listm'.box |> sm'.format
            Fsharp = fun () => chars |> listm'.box |> listm'.to_array' |> sm'.format
            Python = fun () => chars |> listm'.box |> listm'.to_array' |> sm'.format
        }
    if i >= (input |> sm'.length) then
        "parsing.none_of / unexpected end of input / "
        ++# ({ chars' = chars' (); s } |> sm'.format)
        |> Error
    else
        inl ch = input |> sm'.index i
        if chars |> listm'.exists' ((=) ch) |> not
        then Ok (ch, i + 1, s |> update $ch)
        else
            "parsing.none_of / unexpected char / "
            ++# ({ first_char = ch; chars' = chars' (); s } |> sm'.format)
            |> Error

/// ### (<|>)
inl (<|>) forall t. (a : parser t) (b : parser t) : parser t = fun input, i, s =>
    match a (input, i, s) with
    | Ok _ as r => r
    | Error _ => b (input, i, s)

/// ### (|>>)
inl (|>>) p f : parser _ =
    p >> resultm.map fun r, i', s' =>
        f r, i', s'

/// ### many
inl many forall b c. (p : _ * _ * _ -> _ (b * _ * _) c) : parser (list _) = fun input, i0, s0 =>
    // let rec 루프 acc input =
    let rec 루프 (acc : list b) (i : int) (s : parser_state) : result (list b * int * parser_state) string =
        match p (input, i, s) with
        | Ok (x, i', s') =>
            if i' = i
            then "parsing.many / inner parser succeeded without consuming input" |> Error
            else s' |> 루프 (x :: acc) i'
        | Error _ => Ok (acc |> listm.rev, i, s)
    s0 |> 루프 [] i0

/// ### many1_chars
inl many1_chars (p : parser char) : parser string = fun input, i0, s0 =>
    match p (input, i0, s0) with
    | Ok (first, i1, s1) =>
        let rec 루프 (acc : list char) (i : int) (s : parser_state)
            : result (string * int * parser_state) string
            =
            match p (input, i, s) with
            | Ok (c, i', s') =>
                if i' = i
                then "parsing.many1_chars / inner parser succeeded without consuming input" |> Error
                else s' |> 루프 (c :: acc) i'
            | Error _ =>
                Ok (
                    first :: (acc |> listm.rev)
                    |> listm.map sm'.obj_to_string
                    |> listm'.box
                    |> seq.of_list'
                    |> sm'.concat "",
                    i,
                    s
                )
        s1 |> 루프 [] i1
    | Error e => Error e

/// ### many_chars
inl many_chars (p : parser char) : parser string = fun input, i, s =>
    match many1_chars p (input, i, s) with
    | Ok (res, i', s') => Ok (res, i', s')
    | Error _ => Ok ("", i, s)

/// ### many_chars_till
inl many_chars_till (p : parser char) (end_p : parser _) : parser string = fun input, i0, s0 =>
    let rec 루프 (acc : list char) (i : int) (s : parser_state) : result (string * int * parser_state) string =
        inl ok i s =
            Ok (
                acc
                |> listm.rev
                |> listm.map sm'.obj_to_string
                |> listm'.box
                |> seq.of_list'
                |> sm'.concat "",
                i,
                s
            )
        match end_p (input, i, s) with
        | Ok _ => ok i s
        | Error _ =>
            match p (input, i, s) with
            | Ok (_, i', _) when i' = i =>
                "parsing.many_chars_till / inner parser succeeded without consuming input" |> Error
            | Ok (c, i', s') => s' |> 루프 (c :: acc) i'
            | Error _ => ok i s
    s0 |> 루프 [] i0

/// ### many1
inl many1 (p : parser _) : parser (list _) = fun input, i0, s0 =>
    match p (input, i0, s0) with
    | Error e => Error e
    | Ok (first, i1, s1) =>
        let rec 루프 acc (i : int) (s : parser_state) : result (list _ * int * parser_state) string =
            match p (input, i, s) with
            | Ok (x, i', s') =>
                if i' = i
                then "parsing.many1 / inner parser succeeded without consuming input" |> Error
                else s' |> 루프 (x :: acc) i'
            | Error _ => Ok (acc |> listm.rev, i, s)
        s1 |> 루프 [ first ] i1

/// ### many1_strings
inl many1_strings (p : parser _) : parser string = fun input, i, s =>
    match many1 p (input, i, s) with
    | Ok (parts, i', s') =>
        Ok (
            parts
            |> listm.map sm'.obj_to_string
            |> listm'.box
            |> seq.of_list'
            |> sm'.concat "",
            i',
            s'
        )
    | Error e => Error e

/// ### many_strings
inl many_strings (p : parser _) : parser string = fun input, i, s =>
    match many p (input, i, s) with
    | Ok (parts, i', s') =>
        Ok (
            parts
            |> listm.map sm'.obj_to_string
            |> listm'.box
            |> seq.of_list'
            |> sm'.concat "",
            i',
            s'
        )
    | Error _ => Ok ("", i, s)

/// ### choice
inl choice forall t. parsers : parser t = fun input, i, s =>
    let rec 루프 = function
        | [] => "parsing.choice / no parsers succeeded" |> Error
        | (p : _ -> _ (t * int * parser_state) _) :: ps =>
            match p (input, i, s) with
            | Ok _ as r => r
            | Error _ => ps |> 루프
    parsers |> 루프

/// ### between
inl between p_open p_close p_content : parser _ = fun input, i0, s0 =>
    match p_open (input, i0, s0) with
    | Ok (_, i1, s1) =>
        match p_content (input, i1, s1) with
        | Ok (result, i2, s2) =>
            match p_close (input, i2, s2) with
            | Ok (_, i3, s3) => Ok (result, i3, s3)
            | Error e =>
                inl total_len = input |> sm'.length
                inl end1 = (i1 + get_max_context ()) |> min total_len
                inl end2 = (i2 + get_max_context ()) |> min total_len
                inl rest1 = input |> sm'.range (am'.Start i1) (am'.End fun _ => end1)
                inl rest2 = input |> sm'.range (am'.Start i2) (am'.End fun _ => end2)
                "parsing.between / expected closing delimiter / "
                ++# ({ e input rest1 rest2 } |> sm'.format)
                |> Error
        | Error _ => "parsing.between / expected content" |> Error
    | Error e => e |> Error

/// ### sep_by
inl sep_by forall b. p sep : parser (list b) = fun input, i0, s0 =>
    let rec 루프 (acc : list b) (i : int) (s : parser_state) : result (list b * int * parser_state) string =
        match p (input, i, s) with
        | Ok (result, i1, s1) =>
            match sep (input, i1, s1) with
            | Ok (_, i2, s2) => s2 |> 루프 (result :: acc) i2
            | Error _ => Ok ((result :: acc) |> listm.rev, i1, s1)
        | Error _ => Ok (acc |> listm.rev, i, s)
    s0 |> 루프 [] i0

/// ### span_from
inl span_from pred str i0 =
    let rec 루프 (i : int) =
        if i >= (str |> sm'.length)
        then i
        elif pred (str |> sm'.index i)
        then 루프 (i + 1)
        else i
    루프 i0

/// ### spaces1
inl spaces1 () : parser () = fun input, i, s =>
    inl j = i |> span_from ((=) ' ') input
    if j = i
    then "parsing.spaces1 / expected at least one space" |> Error
    else Ok ((), j, s)

/// ### spaces
inl spaces () : parser () = fun input, i, s =>
    Ok ((), i |> span_from ((=) ' ') input, s)

/// ### p_digit
inl p_digit () : parser char = fun input, i, s =>
    if i >= (input |> sm'.length)
    then "parsing.p_digit / unexpected end of input / " ++# ({ s } |> sm'.format) |> Error
    else
        inl c = input |> sm'.index i
        inl cn = c |> try_convert |> optionm'.default_value -1
        if cn >= i32 '0' && cn <= i32 '9'
        then Ok (c, i + 1, s)
        else "parsing.p_digit / unexpected char / " ++# ({ c } |> sm'.format) |> Error

/// ### opt
inl opt p : parser (option _) = fun input, i, s =>
    match p (input, i, s) with
    | Ok (result, i', s') => Ok (result |> Some, i', s')
    | Error _ => Ok (None, i, s)

/// ### rest_of_line
inl rest_of_line () : parser string = fun input, i0, s =>
    inl total_len = input |> sm'.length
    inl j =
        match input |> sm'.index_of_char_from i0 '\n' with
        | -1 => total_len
        | k  => (if k >= i0 then k else i0 + k) |> min total_len
    inl result = input |> sm'.range (am'.Start i0) (am'.End fun _ => j)
    Ok (result, j, s)

/// ### eof
inl eof () : parser () = fun input, i, s =>
    if (input |> sm'.length) = i
    then Ok ((), i, s)
    else
        "parsing.eof / expected end of input / "
        ++# ({ rest = input |> sm'.range (am'.Start i) (am'.End eval) } |> sm'.format)
        |> Error
