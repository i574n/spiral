/// # parsing
open sm'_operators

/// ## fparsec

/// ## parsing

/// ### position

/// ### range
type range =
    {
        from : int
        to : int
    }

type position =
    {
        line : int
        col : int
    }

/// ### parser_state
nominal parser_state =
    {
        line_start : int
        position : position
        input_len : int
    }

/// ### new_parser_state
inl new_parser_state (line_start : i32) (line : i32) (col : i32) (input_len : i32) =
    { line_start position = { line col }; input_len }

/// ### new_parser_state\''
inl new_parser_state' input_len =
    new_parser_state 0 1 1 input_len |> parser_state

/// ### parser
type parser t = string * int * parser_state -> result (t * int * parser_state) string

/// ### slice
inl slice (i0 : int) (i1 : int) (input : string) : string =
    input |> sm'.range (am'.Start i0) (am'.End fun _ => i1)

/// ### parse
inl parse forall t.
    (p : parser t)
    (input : string)
    (s : parser_state)
    : result (t * string * parser_state) string
    =
    p (input, 0, s)
    |> resultm.map fun result, i, s' =>
        result,
        input |> slice i (input |> sm'.length),
        s'

/// ### inc
inl inc (parser_state s) = function
    | '\n' => { line = s.position.line + 1; col = 1 }
    | _ => { s.position with col = s.position.col + 1 }.position

/// ### update_char
inl update_char (parser_state s) (c : char) : parser_state =
    match c with
    | '\n' =>
        { s with
            line_start = s.line_start + s.position.col
            position = { line = s.position.line + 1; col = 1 }
        }
    | _ =>
        { s with
            position = { line = s.position.line; col = s.position.col + 1 }
        }
    |> parser_state

/// ### update
inl update result s =
    inl len = result |> sm'.length
    let rec 루프 (j : int) (parser_state st) =
        if j >= len
        then st |> parser_state
        else
            inl k =
                match result |> sm'.index_of_char_from j '\n' with
                | -1 => -1
                | kk when kk >= j => kk
                | kk => j + kk
            if k = -1 then
                { st with position = { line = st.position.line; col = st.position.col + (len - j) } }
                |> parser_state
            else
                inl st' =
                    if k > j
                    then { st with position = { line = st.position.line; col = st.position.col + (k - j) } }
                    else st
                    |> parser_state
                '\n' |> update_char st' |> 루프 (k + 1)
    s |> 루프 0

/// ### update_span
inl update_span (input : string) (i0 : int) (len : int) (s : parser_state) : parser_state =
    inl endi = i0 + len
    let rec 루프 (j : int) (parser_state st) : parser_state =
        if j >= endi
        then st |> parser_state
        else
            inl k =
                match input |> sm'.index_of_char_from j '\n' with
                | -1 => -1
                | k when k >= j => k
                | k => j + k
            if k = -1 || k >= endi then
                { st with
                    position = { line = st.position.line; col = st.position.col + (endi - j) }
                } |> parser_state
            else
                inl st' =
                    if k <= j
                    then st
                    else
                        { st with
                            position = { line = st.position.line; col = st.position.col + (k - j) }
                        }
                    |> parser_state
                '\n' |> update_char st' |> 루프 (k + 1)
    s |> 루프 i0

/// ### run_parser
inl run_parser parser input =
    input
    |> parse parser
    |> fun parser => parser (new_parser_state' (input |> sm'.length))

/// ### any_char
inl any_char () : parser char = fun input, i, (parser_state st as s) =>
    if i >= st.input_len
    then "parsing.any_char / unexpected end of input / " ++# ({ s } |> sm'.format) |> Error
    else
        inl c = input |> sm'.index i
        Ok (c, i + 1, c |> update_char s)

/// ### get_max_context
inl get_max_context () =
    120

/// ### span_from
inl span_from pred str i0 =
    inl len = str |> sm'.length
    let rec 루프 (i : int) =
        if i >= len
        then i
        elif str |> sm'.index i |> pred
        then 루프 (i + 1)
        else i
    루프 i0

/// ### p_char
inl p_char (c : char) : parser char =
    fun input, i, (parser_state ({ line_start position = { line col } } as st) as s) =>
        if i >= st.input_len
        then "parsing.p_char / unexpected end of input / " ++# ({ c st } |> sm'.format) |> Error
        else
            inl got = input |> sm'.index i
            if got = c
            then Ok (got, i + 1, got |> update_char s)
            else
                inl line_end = i |> span_from ((<>) '\n') input
                inl end = (i + get_max_context ()) |> min line_end
                inl line_slice = input |> slice line_start end
                inl pointer_line = (" " |> sm'.replicate (col - 1)) ++# "^"
                "parsing.p_char / "
                ++# ({ expected = c; line col } |> sm'.format)
                ++# "\n" ++# line_slice
                ++# "\n" ++# pointer_line ++# "\n"
                |> Error

/// ### any_string
inl any_string length : parser string = fun input, i, (parser_state st as s) =>
    if st.input_len - i < length
    then "parsing.any_string / unexpected end of input / " ++# ({ s } |> sm'.format) |> Error
    else Ok (input |> slice i (i + length), i + length, s |> update_span input i length)

/// ### skip_any_string
inl skip_any_string length : parser () = fun input, i, (parser_state st as s) =>
    if st.input_len - i < length
    then "parsing.skip_any_string / unexpected end of input / " ++# ({ s } |> sm'.format) |> Error
    else
        Ok ((), i + length, s |> update_span input i length)

/// ### (>>.)
inl (>>.) forall t u. (a : parser t) (b : parser u) : parser u = fun input, i, s =>
    match a (input, i, s) with
    | Ok (_, i', s') => b (input, i', s')
    | Error e => Error e

/// ### (>>.)
inl (.>>) forall t u. (a : parser t) (b : parser u) : parser t = fun input, i, s =>
    match a (input, i, s) with
    | Ok (ra, i', s') =>
        b (input, i', s')
        |> resultm.map fun _, i'', s'' =>
            ra, i'', s''
    | Error e => Error e

/// ### (.>>.)
inl (.>>.) forall t u. (a : parser t) (b : parser u) : parser (t * u) = fun input, i, s =>
    match a (input, i, s) with
    | Ok (ra, i', s') =>
        b (input,  i', s')
        |> resultm.map fun rb, i'', s'' =>
            (ra, rb), i'', s''
    | Error e => Error e

/// ### (>>%)
inl (>>%) forall t u. (a : parser t) (b : u) : parser u =
    a >> resultm.map fun _, i', s' =>
        b, i', s'

/// ### none_of
inl none_of (chars : list char) : parser char = fun input, i, (parser_state st as s) =>
    inl chars' () =
        chars |> listm'.box |> listm'.to_array' |> sm'.format
    if i >= st.input_len
    then "parsing.none_of / unexpected end of input / " ++# ({ chars' = chars' (); s } |> sm'.format) |> Error
    else
        inl ch = input |> sm'.index i
        if chars |> listm'.exists' ((=) ch) |> not
        then Ok (ch, i + 1, ch |> update_char s)
        else
            "parsing.none_of / unexpected char / "
            ++# ({ first_char = ch; chars' = chars' (); s } |> sm'.format)
            |> Error

/// ### (<|>)
inl (<|>) forall t. (a : parser t) (b : parser t) : parser t = fun input, i, s =>
    match a (input, i, s) with
    | Ok _ as r => r
    | Error _ => b (input, i, s)

/// ### (|>>)
inl (|>>) p f : parser _ =
    p >> resultm.map fun r, i', s' =>
        f r, i', s'

/// ### many
inl many forall b c.
    (p : _ * _ * _ -> _ (b * _ * _) c)
    : parser (list _)
    =
    fun input, i0, (parser_state st as s0) =>
        let rec 루프 (acc : list b) (i : int) (fuel : int) (s : parser_state)
            : result (list b * int * parser_state) string
            =
            if fuel <= 0
            then "parsing.many / out of fuel (probable zero-length loop)" |> Error
            else
                match p (input, i, s) with
                | Ok (x, i', s') when i' = i =>
                    "parsing.many / inner parser succeeded without consuming input" |> Error
                | Ok (x, i', s') => s' |> 루프 (x :: acc) i' (fuel - 1)
                | Error _ => Ok (acc |> listm.rev, i, s)
        s0 |> 루프 [] i0 (st.input_len - i0 + 2)

/// ### many1_chars
inl many1_chars (p : parser char) : parser string = fun input, i0, s0 =>
    match p (input, i0, s0) with
    | Error e => Error e
    | Ok (_, i1, s1) =>
        let rec 루프 (i : int) (s : parser_state) : result (string * int * parser_state) string =
            match p (input, i, s) with
            | Ok (_, i', s') =>
                if i' = i
                then "parsing.many1_chars / inner parser succeeded without consuming input" |> Error
                else s' |> 루프 i'
            | Error _ => Ok (input |> slice i0 i, i, s)
        s1 |> 루프 i1

/// ### many_chars
inl many_chars (p : parser char) : parser string = fun input, i, s =>
    match many1_chars p (input, i, s) with
    | Ok (res, i', s') => Ok (res, i', s')
    | Error _ => Ok ("", i, s)

/// ### many_chars_till
inl many_chars_till (p : parser char) (end_p : parser _) : parser string = fun input, i0, s0 =>
    let rec 루프 (i : int) (s : parser_state) : result (string * int * parser_state) string =
        match end_p (input, i, s) with
        | Ok _ => Ok ((if i > i0 then input |> slice i0 i else ""), i, s)
        | Error _ =>
            match p (input, i, s) with
            | Ok (_, i', s') =>
                if i' = i
                then "parsing.many_chars_till / inner parser succeeded without consuming input" |> Error
                else s' |> 루프 i'
            | Error _ => Ok ((if i > i0 then input |> slice i0 i else ""), i, s)
    s0 |> 루프 i0

/// ### many1
inl many1 (p : parser _) : parser (list _) = fun input, i0, (parser_state st as s0) =>
    match p (input, i0, s0) with
    | Error e => e |> Error
    | Ok (first, i1, s1) =>
        inl fuel_max = st.input_len - i1 + 2
        let rec 루프 acc (i : int) (fuel : int) s : result (list _ * int * parser_state) string =
            if fuel <= 0
            then "parsing.many1 / out of fuel (probable zero-length loop)" |> Error
            else
                match p (input, i, s) with
                | Ok (x, i', s') =>
                    if i' = i
                    then "parsing.many1 / inner parser succeeded without consuming input" |> Error
                    else s' |> 루프 (x :: acc) i' (fuel - 1)
                | Error _ => Ok (acc |> listm.rev, i, s)
        s1 |> 루프 [ first ] i1 fuel_max

/// ### many1_strings
inl many1_strings (p : parser _) : parser string = fun input, i0, (parser_state st as s0) =>
    match p (input, i0, s0) with
    | Error e => e |> Error
    | Ok (r0, i1, s1) =>
        inl fuel_max = st.input_len - i1 + 2
        let rec 루프 (acc : list string) (i : int) (fuel : int) s : result (string * int * _) string =
            if fuel <= 0
            then "parsing.many1_strings / out of fuel (probable zero-length loop)" |> Error
            else
                match p (input, i, s) with
                | Error _ => Ok (acc |> listm.rev |> sm'.concat_list "", i, s)
                | Ok (r, i', s') =>
                    if i' = i
                    then "parsing.many1_strings / inner parser succeeded without consuming input" |> Error
                    else s' |> 루프 ($r :: acc) i' (fuel - 1)
        s1 |> 루프 [ $r0 ] i1 fuel_max

/// ### many_strings
inl many_strings (p : parser _) : parser string = fun input, i0, (parser_state st as s0) =>
    match p (input, i0, s0) with
    | Error _ => Ok ("", i0, s0)
    | Ok (r0, i1, s1) when i1 = i0 => "parsing.many_strings / first inner parser consumed no input" |> Error
    | Ok (r0, i1, s1) =>
        inl fuel_max = st.input_len - i1 + 2
        let rec 루프 (acc : list string) (i : int) (fuel : int) s : result (string * int * _) string =
            if fuel <= 0
            then "parsing.many_strings / out of fuel (probable zero-length loop)" |> Error
            else
                match p (input, i, s) with
                | Ok (r, i', s') when i' = i =>
                    "parsing.many_strings / inner parser succeeded without consuming input" |> Error
                | Ok (r, i', s') => s' |> 루프 ($r :: acc) i' (fuel - 1)
                | Error _ => Ok ($r0 :: (acc |> listm.rev) |> sm'.concat_list "", i, s)
        s1 |> 루프 [] i1 fuel_max

/// ### choice
inl choice forall t. parsers : parser t = fun input, i, s =>
    let rec 루프 = function
        | [] => "parsing.choice / no parsers succeeded" |> Error
        | (p : _ -> _ (t * int * parser_state) _) :: ps =>
            match p (input, i, s) with
            | Ok _ as r => r
            | Error _ => ps |> 루프
    parsers |> 루프

/// ### between
inl between p_open p_close p_content : parser _ = fun input, i0, s0 =>
    match p_open (input, i0, s0) with
    | Ok (_, i1, s1) =>
        match p_content (input, i1, s1) with
        | Ok (result, i2, s2) =>
            match p_close (input, i2, s2) with
            | Ok (_, i3, s3) => Ok (result, i3, s3)
            | Error e =>
                inl total_len = input |> sm'.length
                inl end1 = (i1 + get_max_context ()) |> min total_len
                inl end2 = (i2 + get_max_context ()) |> min total_len
                inl rest1 = input |> slice i1 end1
                inl rest2 = input |> slice i2 end2
                "parsing.between / expected closing delimiter / "
                ++# ({ e input rest1 rest2 } |> sm'.format)
                |> Error
        | Error _ =>
            match p_close (input, i1, s1) with
            | Ok (_, i3, s3) => Ok ("", i3, s3)
            | Error _ =>
                inl total_len = input |> sm'.length
                inl end1 = (i1 + get_max_context ()) |> min total_len
                inl rest1 = input |> slice i1 end1
                "parsing.between / expected content or closing delimiter / "
                ++# ({ rest1 } |> sm'.format)
                |> Error
    | Error e => e |> Error

/// ### sep_by
inl sep_by forall b. p sep : parser (list b) = fun input, i0, s0 =>
    match p (input, i0, s0) with
    | Error _ => Ok ([], i0, s0)
    | Ok (first, i1, s1) =>
        let rec 루프 (acc : list b) (i : int) s : result (list b * int * parser_state) string =
            match sep (input, i, s) with
            | Ok (_, j, s') =>
                if j = i
                then "parsing.sep_by / separator consumed no input" |> Error
                else
                    match p (input, j, s') with
                    | Ok (x, k, s'') => s'' |> 루프 (x :: acc) k
                    | Error _ => Ok (acc |> listm.rev, i, s)
            | Error _ => Ok (acc |> listm.rev, i, s)
        s1 |> 루프 [ first ] i1

/// ### is_space
inl is_space c =
    c = ' ' || c = '\t' || c = '\r'

/// ### spaces1
inl spaces1 () : parser () = fun input, i, s =>
    inl j = i |> span_from is_space input
    if j = i
    then "parsing.spaces1 / expected at least one space" |> Error
    else Ok ((), j, s |> update_span input i (j - i))

/// ### spaces
inl spaces () : parser () = fun input, i, s =>
    inl j = i |> span_from is_space input
    Ok ((), j, s |> update_span input i (j - i))

/// ### p_digit
inl p_digit () : parser char = fun input, i, (parser_state st as s) =>
    if i >= st.input_len
    then "parsing.p_digit / unexpected end of input / " ++# ({ s } |> sm'.format) |> Error
    else
        match input |> sm'.index i with
        | '0' | '1' | '2' | '3' | '4' | '5' | '6' | '7' | '8' | '9' as c => Ok (c, i + 1, c |> update_char s)
        | c => "parsing.p_digit / unexpected char / " ++# ({ c } |> sm'.format) |> Error

/// ### opt
inl opt p : parser (option _) = fun input, i, s =>
    match p (input, i, s) with
    | Ok (result, i', s') => Ok (result |> Some, i', s')
    | Error _ => Ok (None, i, s)

/// ### rest_of_line
inl rest_of_line () : parser string = fun input, i0, (parser_state st as s) =>
    inl j =
        match input |> sm'.index_of_char_from i0 '\n' with
        | -1 => st.input_len
        | k => if k >= i0 then k else i0 + k
    Ok (input |> slice i0 j, j, s |> update_span input i0 (j - i0))

/// ### eof
inl eof () : parser () = fun input, i, (parser_state st as s) =>
    if st.input_len = i
    then Ok ((), i, s)
    else
        "parsing.eof / expected end of input / "
        ++# ({ rest = input |> slice i st.input_len } |> sm'.format)
        |> Error
