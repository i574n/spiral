/// # parsing
open sm'_operators

/// ## fparsec

/// ## parsing

/// ### position

/// ### range
type range =
    {
        from : int
        to : int
    }

type position =
    {
        line : int
        col : int
    }

/// ### parser_state
nominal parser_state =
    {
        line_start : int
        position : position
        text_length : int
    }

/// ### new_parser_state
inl new_parser_state (line_start : i32) (line : i32) (col : i32) (text_length : i32) =
    { line_start position = { line col }; text_length }

/// ### new_parser_state\''
inl new_parser_state' text_length =
    new_parser_state 0 1 1 text_length |> parser_state

/// ### parser
type parser t = string * int * parser_state -> result ((() -> t) * int * parser_state) (() -> string)

/// ### slice
inl slice (start : int) (end : int) (t : string) : string =
    t
    |> sm'.range (am'.Start start) (am'.End fun _ => end)
    |> trace_format Verbose fun r =>
        "parsing.slice", { start end t_len = ##t; r_length = ##r }

/// ### parse
inl parse forall t.
    (p : parser t)
    (t : string)
    (s : parser_state)
    : result ((() -> t) * (() -> string) * parser_state) (() -> string)
    =
    p (t, 0, s)
    |> resultm.map fun result, i, (parser_state s' as s) =>
        result,
        (fun () => t |> slice i s'.text_length),
        s

/// ### update_char
inl update_char (parser_state s) (c : char) : parser_state =
    match c with
    | '\n' =>
        { s with
            line_start = s.line_start + s.position.col
            position = { line = s.position.line + 1; col = 1 }
        }
    | _ =>
        { s with
            position = { line = s.position.line; col = s.position.col + 1 }
        }
    |> parser_state
    |> trace_format Verbose fun r => "parsing.update_char", { c s r }

/// ### update_span
inl update_span (t : string) (i : int) (len : int) (parser_state s' as s) : parser_state =
    inl endi = i + len
    let rec 루프 (i' : int) (last_nl : int) (count : int) =
        trace Verbose
            (fun () => "parsing.update_span / 루프")
            (fun () => { i len endi i' last_nl count t_len = ##t; s })
        if i' >= endi
        then last_nl, count
        else
            match t |> sm'.index i' with
            | '\n' => 루프 (i' + 1) i' (count + 1)
            | _ => 루프 (i' + 1) last_nl count
    inl last_nl, n = 루프 i -1 0
    if n = 0
    then { s' with position = { line = s'.position.line; col = s'.position.col + len } }
    else
        { s' with
            line_start = last_nl + 1
            position =
                {
                    line = s'.position.line + n
                    col = endi - last_nl
                }
            text_length = s'.text_length
        }
    |> parser_state
    |> trace_format Verbose fun r =>
        "parsing.update_span", { i len endi last_nl n t_len = ##t; s r }

/// ### update
inl update t s =
    s
    |> update_span t 0 ##t
    |> trace_format Verbose fun r => "parsing.update", { t s r }

/// ### advance_while
inl advance_while (fn : char -> bool) (t : string) (i : int) (parser_state s' as s)
    : int * parser_state
    =
    if i >= s'.text_length
    then i, s
    else
        inl i' = i |> sm'.span_from fn t
        inl i' =
            if i' > s'.text_length
            then s'.text_length
            else i'
        inl consumed = i' - i
        if consumed = 0
        then i, s
        else i', s |> update_span t i consumed
    |> trace_format Verbose fun r =>
        "parsing.advance_while", { i t_len = ##t; s r }

/// ### run_parser
inl run_parser p t =
    t
    |> parse p
    |> fun run => ##t |> new_parser_state' |> run
    |> resultm.map fun a, b, s => a (), b (), s

/// ### any_char
inl any_char () : parser char = fun t, i, (parser_state s' as s) =>
    if i >= s'.text_length then
        fun () => "parsing.any_char / unexpected end of t / " ++#? { s }
        |> Error
    else
        inl c = t |> sm'.index i
        trace Verbose (fun () => "parsing.any_char") (fun () => { c s })
        Ok ((fun () => c), i + 1, c |> update_char s)
    |> trace_format Verbose fun r => "parsing.any_char", { i t_len = ##t; s r }

/// ### get_max_context
inl get_max_context () =
    80

/// ### p_char
inl p_char (c : char) : parser char =
    fun t, i, (parser_state ({ line_start position = { line col } } as s') as s) =>
        trace Verbose (fun () => "parsing.p_char") (fun () => { c t_len = ##t; i s })
        if i >= s'.text_length then
            fun () => "parsing.p_char / unexpected end of text / " ++#? { c s' }
            |> Error
        else
            inl got = t |> sm'.index i
            if got = c
            then Ok ((fun () => got), i + 1, got |> update_char s)
            else
                fun () =>
                    inl line_end = i |> sm'.span_from ((<>) '\n') t
                    inl end = (i + get_max_context ()) |> min line_end
                    inl line_slice = t |> slice line_start end
                    inl new_line =
                        inl len = ##line_slice
                        if len > 0 && (line_slice |> sm'.index (len - 1)) = '\n' then "" else "\n"
                    inl pointer_line = (" " |> sm'.replicate (col - 1)) ++# "^"
                    "parsing.p_char / "
                    ++#? { expected = c; line col }
                    ++# "\n" ++# line_slice
                    ++# new_line
                    ++# pointer_line ++# "\n"
                |> Error

/// ### any_string
inl any_string len : parser string = fun t, i, (parser_state s' as s) =>
    trace Verbose (fun () => "parsing.any_string") (fun () => { t_len = ##t; i s })
    if s'.text_length - i >= len
    then Ok ((fun () => t |> slice i (i + len)), i + len, s |> update_span t i len)
    else
        fun () => "parsing.any_string / unexpected end of text / " ++#? { s }
        |> Error

/// ### skip_any_string
inl skip_any_string len : parser () = fun t, i, (parser_state s' as s) =>
    trace Verbose (fun () => "parsing.skip_any_string") (fun () => { t_len = ##t; i s })
    if s'.text_length - i >= len
    then Ok (id, i + len, s |> update_span t i len)
    else
        fun () => "parsing.skip_any_string / unexpected end of text / " ++#? { s }
        |> Error

/// ### skip_many
inl skip_many forall t. (p : parser t) : parser () = fun t, i, s =>
    trace Verbose (fun () => "parsing.skip_many") (fun () => { t_len = ##t; i s })
    let rec 루프 (i' : int) (s' : parser_state) =
        trace Verbose
            fun () => "parsing.skip_many / 루프"
            fun () => { t_len = ##t; i s i' s' }
        match p (t, i', s') with
        | Error _ => Ok (id : () -> (), i', s')
        | Ok (_, i'', s'') =>
            if i'' <> i'
            then s'' |> 루프 i''
            else
                fun () => "parsing.skip_many / inner parser consumed no text"
                |> Error
    s |> 루프 i

/// ### skip_many1
inl skip_many1 forall t. (a : parser t) : parser () = fun t, i, s =>
    trace Verbose (fun () => "parsing.skip_many1") (fun () => { t_len = ##t; i s })
    match a (t, i, s) with
    | Error e => e |> Error
    | Ok (_, i', s') =>
        if i' <> i
        then skip_many a (t, i', s')
        else
            fun () => "parsing.skip_many1 / inner parser consumed no text"
            |> Error

/// ### (>>.)
inl (>>.) forall t u. (a : parser t) (b : parser u) : parser u = fun t, i, s =>
    trace Verbose (fun () => "parsing.(>>.)") (fun () => { t_len = ##t })
    match a (t, i, s) with
    | Ok (_, i', s') => b (t, i', s')
    | Error e => e |> Error

/// ### (.>>)
inl (.>>) forall t u. (a : parser t) (b : parser u) : parser t = fun t, i, s =>
    trace Verbose (fun () => "parsing.(.>>)") (fun () => { t_len = ##t })
    match a (t, i, s) with
    | Error e => e |> Error
    | Ok (ra, i', s') =>
        b (t, i', s')
        |> resultm.map fun _, i'', s'' =>
            ra, i'', s''

/// ### (.>>.)
inl (.>>.) forall t u. (a : parser t) (b : parser u) : parser ((() -> t) * (() -> u)) = fun t, i, s =>
    trace Verbose (fun () => "parsing.(.>>.)") (fun () => { t_len = ##t })
    match a (t, i, s) with
    | Error e => e |> Error
    | Ok (ra, i', s') =>
        b (t, i', s')
        |> resultm.map fun rb, i'', s'' =>
            (fun () => ra, rb), i'', s''

/// ### (>>%)
inl (>>%) forall t u. (a : parser t) (b : u) : parser u =
    trace Verbose (fun () => "parsing.(>>%)") (fun () => { b })
    a >> resultm.map fun _, i', s' =>
        (fun () => b), i', s'

/// ### none_of
inl none_of (chars : list char) : parser char = fun t, i, (parser_state s' as s) =>
    trace Verbose (fun () => "parsing.none_of") (fun () => { chars t_len = ##t; i s })
    inl chars' () =
        chars |> listm'.box |> listm'.to_array' |> sm'.format
    if i >= s'.text_length then
        fun () => "parsing.none_of / unexpected end of text / " ++#? { chars' = chars' (); s }
        |> Error
    else
        inl ch = t |> sm'.index i
        if chars |> listm'.exists' ((=) ch) |> not
        then Ok ((fun () => ch), i + 1, ch |> update_char s)
        else
            fun () =>
                "parsing.none_of / unexpected char / "
                ++#? { first_char = ch; chars' = chars' (); s }
            |> Error

/// ### (<|>)
inl (<|>) forall t. (a : parser t) (b : parser t) : parser t = fun t, i, s =>
    trace Verbose (fun () => "parsing.(<|>)") (fun () => { t_len = ##t; i s })
    match a (t, i, s) with
    | Ok _ as r => r
    | Error _ => b (t, i, s)

/// ### (|>>)
inl (|>>) p f : parser _ =
    trace Verbose (fun () => "parsing.(|>>)") (fun () => {})
    p >> resultm.map fun r, i', s' =>
        f r, i', s'

/// ### many
inl many forall b c.
    (p : _ * _ * _ -> _ ((() -> b) * _ * _) c)
    : parser (list _)
    =
    fun t, i, s =>
        trace Verbose (fun () => "parsing.many") (fun () => { t_len = ##t })
        let rec 루프 (acc : list b) (i' : int) (s' : parser_state)
            : result ((() -> list b) * int * parser_state) _
            =
            trace Verbose
                fun () => "parsing.many / 루프"
                fun () => { t_len = ##t; i' s' }
            match p (t, i', s') with
            | Error _ => Ok ((fun () => acc |> listm.rev), i', s')
            | Ok (x, i'', s'') when i'' > i' => s'' |> 루프 (x () :: acc) i''
            | Ok _ =>
                fun () => "parsing.many / inner parser succeeded without consuming text"
                |> Error
        s |> 루프 [] i

/// ### many1_chars
inl many1_chars (p : parser char) : parser string = fun t, i, s =>
    trace Verbose (fun () => "parsing.many1_chars") (fun () => { t_len = ##t; i s })
    match p (t, i, s) with
    | Error e => e |> Error
    | Ok (_, i', s') =>
        let rec 루프 (i'' : int) (s'' : parser_state) : result ((() -> string) * int * parser_state) _ =
            trace Verbose
                fun () => "parsing.many1_chars / 루프"
                fun () => { t_len = ##t; i s i'' s'' }
            match p (t, i'', s'') with
            | Error _ => Ok ((fun () => t |> slice i i''), i'', s'')
            | Ok (_, i''', s''') =>
                if i''' <> i''
                then s''' |> 루프 i'''
                else
                    fun () => "parsing.many1_chars / inner parser succeeded without consuming text"
                    |> Error
        s' |> 루프 i'

/// ### many_chars
inl many_chars (p : parser char) : parser string = fun t, i, s =>
    trace Verbose (fun () => "parsing.many_chars") (fun () => { t_len = ##t; i s })
    match many1_chars p (t, i, s) with
    | Ok (res, i', s') => Ok (res, i', s')
    | Error _ => Ok ((fun () => ""), i, s)

/// ### many_chars_till
inl many_chars_till (p : parser char) (end_p : parser _) = fun t, i, (parser_state s' as s) =>
    trace Verbose (fun () => "parsing.many_chars_till") (fun () => { t_len = ##t; i s })
    let rec 루프 (i' : int) (s'' : parser_state) : result ((() -> string) * int * parser_state) (() -> string) =
        trace Verbose
            fun () => "parsing.many_chars_till"
            fun () => { t_len = ##t; i s i' s'' }
        if i' >= s'.text_length
        then Ok ((fun () => if i' > i then t |> slice i i' else ""), i', s'')
        else
            inl i'', s''' = s'' |> advance_while (fun c => c <> '\n') t i'
            if i'' >= s'.text_length
            then Ok ((fun () => if i'' > i then t |> slice i i'' else ""), i'', s''')
            else
                match end_p (t, i'', s''') with
                | Ok _ => Ok ((fun () => if i'' > i then t |> slice i i'' else ""), i'', s''')
                | Error _ =>
                    match p (t, i'', s''') with
                    | Error _ => Ok ((fun () => if i'' > i then t |> slice i i'' else ""), i'', s''')
                    | Ok (_, i''', s'''') when i''' > i'' => s'''' |> 루프 i'''
                    | Ok _ =>
                        fun () => "parsing.many_chars_till / inner parser succeeded without consuming text"
                        |> Error
    s |> 루프 i

/// ### many1
inl many1 (p : parser _) : parser (list _) = fun t, i, s =>
    trace Verbose (fun () => "parsing.many1") (fun () => { t_len = ##t; i s })
    match p (t, i, s) with
    | Error e => e |> Error
    | Ok (first, i', s') =>
        let rec 루프 acc (i'' : int) s'' : result ((() -> list _) * int * parser_state) _ =
            trace Verbose
                fun () => "parsing.many1 / 루프"
                fun () => { t_len = ##t; i s i'' s'' }
            match p (t, i'', s'') with
            | Error _ => Ok ((fun () => acc |> listm.rev), i'', s'')
            | Ok (x, i''', s''') when i''' > i'' => s''' |> 루프 (x () :: acc) i'''
            | Ok _ =>
                fun () => "parsing.many1 / inner parser succeeded without consuming text"
                |> Error
        s' |> 루프 [ first () ] i'

/// ### many1_strings
inl many1_strings (p : parser _) : parser string = fun t, i, s =>
    trace Verbose (fun () => "parsing.many1_strings") (fun () => { t_len = ##t })
    match p (t, i, s) with
    | Error e => e |> Error
    | Ok (r, i', s') =>
        let rec 루프 (acc : list string) (i'' : int) s'' : result ((() -> string) * int * _) _ =
            trace Verbose
                fun () => "parsing.many1_strings / 루프"
                fun () => { t_len = ##t; i'' s'' }
            match p (t, i'', s'') with
            | Error _ => Ok ((fun () => acc |> listm.rev |> sm'.concat_list ""), i'', s'')
            | Ok (r', i''', s''') when i''' > i => s''' |> 루프 (#?(r' ()) :: acc) i'''
            | Ok _ =>
                fun () => "parsing.many1_strings / inner parser succeeded without consuming text"
                |> Error
        s' |> 루프 [ #?(r ()) ] i'

/// ### many_strings
inl many_strings (p : parser _) : parser string = fun t, i, s =>
    trace Verbose (fun () => "parsing.many_strings") (fun () => { t_len = ##t })
    match p (t, i, s) with
    | Error _ => Ok ((fun () => ""), i, s)
    | Ok (_, i', _) when i' = i =>
        fun () => "parsing.many_strings / first inner parser consumed no text"
        |> Error
    | Ok (r, i', s') =>
        let rec 루프 (acc : list string) (i' : int) s' : result ((() -> string) * int * _) _ =
            trace Verbose
                fun () => "parsing.many_strings / 루프"
                fun () => { t_len = ##t; i' s' }
            match p (t, i', s') with
            | Error _ => Ok ((fun () => #?(r ()) :: (acc |> listm.rev) |> sm'.concat_list ""), i', s')
            | Ok (r', i'', s'') when i'' > i' => s'' |> 루프 (#?(r' ()) :: acc) i''
            | Ok _ =>
                fun () => "parsing.many_strings / inner parser succeeded without consuming text"
                |> Error
        s' |> 루프 [] i'

/// ### choice
inl choice forall t. ps : parser t = fun t, i, s =>
    trace Verbose
        (fun () => "parsing.choice")
        (fun () => { t_len = ##t; i s ps_length = ps |> listm.length : int })
    let rec 루프 = function
        | [] =>
            fun () => "parsing.choice / no parsers succeeded"
            |> Error
        | (p : _ -> _ ((() -> t) * int * parser_state) _) :: ps' =>
            trace Verbose
                (fun () => "parsing.choice / 루프")
                (fun () => { t_len = ##t; i s ps'_length = ps' |> listm.length : int })
            match p (t, i, s) with
            | Ok _ as r => r
            | Error _ => ps' |> 루프
    ps |> 루프

/// ### between
inl between p_open p_close p_content : parser _ = fun t, i, s =>
    trace Verbose (fun () => "parsing.between") (fun () => { t_len = ##t; i s })
    match p_open (t, i, s) with
    | Ok (_, i', s') =>
        match p_content (t, i', s') with
        | Ok (result, i'', s'') =>
            match p_close (t, i'', s'') with
            | Ok (_, i''', s''') => Ok (result, i''', s''')
            | Error e =>
                fun () =>
                    inl t_len = ##t
                    inl end' = (i' + get_max_context ()) |> min t_len
                    inl end'' = (i'' + get_max_context ()) |> min t_len
                    inl rest' = t |> slice i' end'
                    inl rest'' = t |> slice i'' end''
                    "parsing.between / expected closing delimiter / " ++#? { e t rest' rest'' }
                |> Error
        | Error _ =>
            match p_close (t, i', s') with
            | Ok (_, i''', s''') => Ok ((fun () => ""), i''', s''')
            | Error _ =>
                fun () =>
                    inl end' = (i' + get_max_context ()) |> min ##t
                    inl rest' = t |> slice i' end'
                    "parsing.between / expected content or closing delimiter / " ++#? { rest' }
                |> Error
    | Error e => e |> Error

/// ### sep_by
inl sep_by forall b. p sep : parser (list b) = fun t, i, s =>
    trace Verbose (fun () => "parsing.sep_by") (fun () => { t_len = ##t; i s })
    match p (t, i, s) with
    | Error _ => Ok ((fun () => []), i, s)
    | Ok (first, i', s') =>
        let rec 루프 (acc : list b) (i'' : int) s'' : result ((() -> list b) * int * parser_state) _ =
            trace Verbose
                (fun () => "parsing.sep_by / 루프")
                (fun () => { t_len = ##t; i s i'' s'' })
            match sep (t, i'', s'') with
            | Error _ => Ok ((fun () => acc |> listm.rev), i'', s'')
            | Ok (_, i''', s''') =>
                if i''' = i'' then
                    fun () => "parsing.sep_by / separator consumed no text"
                    |> Error
                else
                    match p (t, i''', s''') with
                    | Ok (x, i'''', s'''') => s'''' |> 루프 (x () :: acc) i''''
                    | Error _ => Ok ((fun () => acc |> listm.rev), i'', s'')
        s' |> 루프 [ first () ] i'

/// ### sep_end_by
inl sep_end_by forall b. p sep : parser (list b) = fun t, i, s =>
    trace Verbose (fun () => "parsing.sep_end_by") (fun () => { t_len = ##t; i s })
    let rec 루프 acc i' s' =
        trace Verbose
            (fun () => "parsing.sep_end_by / 루프")
            (fun () => { t_len = ##t; i s i' s' })
        match p (t, i', s') with
        | Error _ => Ok ((fun () => acc |> listm.rev), i', s')
        | Ok (x, i'', s'') =>
            if i'' = i' then
                fun () => "parsing.sep_end_by / element parser consumed no text"
                |> Error
            else
                inl acc' = x () :: acc
                match sep (t, i'', s'') with
                | Error _ => Ok ((fun () => acc' |> listm.rev), i'', s'')
                | Ok (_, i''', s''') =>
                    if i''' <> i''
                    then s''' |> 루프 acc' i'''
                    else
                        fun () => "parsing.sep_end_by / separator consumed no text"
                        |> Error
    s |> 루프 [] i

/// ### is_space
inl is_space c =
    c = ' ' || c = '\t' || c = '\r'

/// ### spaces1
inl spaces1 () : parser () = fun t, i, (parser_state s' as s) =>
    inl i', s' = s |> advance_while is_space t i
    trace Verbose (fun () => "parsing.spaces1") (fun () => { t_len = ##t; i s i' s' })
    if i' <> i
    then Ok (id, i', s')
    else
        fun () =>
            inl preview_end = (i + get_max_context ()) |> min s'.text_length
            "parsing.spaces1 / expected at least one space / "
            ++#? { rest = t |> slice i preview_end }
        |> Error

/// ### spaces
inl spaces () : parser () = fun t, i, s =>
    inl i', s' = s |> advance_while is_space t i
    trace Verbose (fun () => "parsing.spaces") (fun () => { t_len = ##t; i i' s s' })
    Ok (id, i', s')

/// ### p_digit
inl p_digit () : parser char = fun t, i, (parser_state s' as s) =>
    trace Verbose (fun () => "parsing.p_digit") (fun () => { t_len = ##t; i s })
    if i >= s'.text_length then
        fun () => "parsing.p_digit / unexpected end of text / " ++#? { s }
        |> Error
    else
        match t |> sm'.index i with
        | '0' | '1' | '2' | '3' | '4' | '5' | '6' | '7' | '8' | '9' as c =>
            Ok ((fun () => c), i + 1, c |> update_char s)
        | c =>
            fun () => "parsing.p_digit / unexpected char / " ++#? { c }
            |> Error

/// ### opt
inl opt p : parser (option _) = fun t, i, s =>
    trace Verbose (fun () => "parsing.opt") (fun () => { t_len = ##t })
    match p (t, i, s) with
    | Ok (r, i', s') => Ok ((fun () => r |> Some), i', s')
    | Error _ => Ok ((fun () => None), i, s)

/// ### rest_of_line
inl rest_of_line () : parser string = fun t, i, s =>
    trace Verbose (fun () => "parsing.rest_of_line") (fun () => { t_len = ##t })
    inl i'', s' = s |> advance_while ((<>) '\n') t i
    Ok ((fun () => t |> slice i i''), i'', s')

/// ### eof
inl eof () : parser () = fun t, i, (parser_state s' as s) =>
    trace Verbose (fun () => "parsing.eof") (fun () => { t_len = ##t })
    if s'.text_length = i
    then Ok (id, i, s)
    else
        fun () =>
            "parsing.eof / expected end of text / "
            ++#? { rest = t |> slice i s'.text_length }
        |> Error

/// ### p_string
inl p_string (str : string) : parser string = fun t, i, (parser_state s' as s) =>
    trace Verbose (fun () => "parsing.p_string") (fun () => { t_len = ##t })
    inl len = ##str
    if s'.text_length - i < len then
        fun () => "parsing.p_string / unexpected end of text / " ++#? { expected = str; s }
        |> Error
    else
        let rec eq k =
            if k >= len
            then true
            else t |> sm'.index (i + k) = str |> sm'.index k && eq (k + 1)
        if eq 0
        then Ok ((fun () => t |> slice i (i + len)), i + len, s |> update_span t i len)
        else
            fun () =>
                inl preview_end = (i + get_max_context ()) |> min s'.text_length
                inl rest = t |> slice i preview_end
                inl got = t |> slice i (i + len)
                "parsing.p_string / unexpected string / "
                ++#? { expected = str; got rest s }
            |> Error

/// ### new_line
inl new_line () : parser char = fun t, i, (parser_state s' as s) =>
    trace Verbose (fun () => "parsing.new_line") (fun () => { t_len = ##t })
    if i >= s'.text_length then
        fun () => "parsing.new_line / unexpected end of text / " ++#? { s }
        |> Error
    else
        inl c = t |> sm'.index i
        if c = '\n'
        then Ok ((fun () => c), i + 1, c |> update_char s)
        else
            fun () =>
                inl preview_end = (i + get_max_context ()) |> min s'.text_length
                inl rest = t |> slice i preview_end
                "parsing.new_line / expected new line char / "
                ++#? { first_char = c; rest s }
            |> Error

/// ### many_till
inl many_till forall b c. (p : parser b) (end_p : parser c) : parser _ = fun t, i, s =>
    trace Verbose (fun () => "parsing.many_till") (fun () => { i t_len = ##t })
    let rec 루프 (acc : list b) (i' : int) s' : result (_ * int * parser_state) _ =
        trace Verbose
            (fun () => "parsing.many_till / loop")
            (fun () => { i' acc_len = acc |> listm.length : int })
        match end_p (t, i', s') with
        | Ok (_, i'', s'') => Ok ((fun () => acc |> listm.rev), i'', s'')
        | Error _ =>
            match p (t, i', s') with
            | Ok (x, i'', s'') =>
                if i'' <> i'
                then s'' |> 루프 (x () :: acc) i''
                else
                    fun () => "parsing.many_till / inner parser succeeded without consuming text"
                    |> Error
            | Error e => e |> Error
    s |> 루프 [] i

/// ### p_return
inl p_return forall t. (x : t) : parser t = fun t, i, s =>
    trace Verbose (fun () => "parsing.p_return") (fun () => { t_len = ##t })
    Ok ((fun () => x), i, s)

/// ### attempt
inl attempt forall t. (p : parser t) : parser t = fun t, i, s =>
    trace Verbose (fun () => "parsing.attempt") (fun () => { t_len = ##t })
    match p (t, i, s) with
    | Ok (r, i', s') => Ok (r, i', s')
    | Error e => e |> Error

/// ### look_ahead
inl look_ahead (p : parser _) : parser _ = fun t, i, s =>
    trace Verbose (fun () => "parsing.look_ahead") (fun () => { t_len = ##t })
    match p (t, i, s) with
    | Ok (x, _, _) => Ok (x, i, s)
    | Error e => e |> Error
    |> trace_format Verbose fun r => "parsing.look_ahead", { t_len = ##t; r}

/// ### pipe2
inl pipe2 forall a b c. (p1 : parser a) (p2 : parser b) (f : ((() -> a) * (() -> b)) -> c) : parser c =
    p1 .>>. p2 |>> fun r => fun () =>
        trace Verbose (fun () => "parsing.pipe2") (fun () => {})
        r () |> f

/// ### new_lines
inl new_lines () : parser () = fun t, i, s =>
    trace Verbose (fun () => "parsing.new_lines") (fun () => { t_len = ##t })
    inl i', s' = s |> advance_while ((=) '\n') t i
    Ok (id, i', s')
    |> trace_format Verbose fun r => "parsing.new_lines", { t_len = ##t; r}

/// ### new_lines1
inl new_lines1 () : parser () = fun t, i, (parser_state s' as s) =>
    trace Verbose (fun () => "parsing.new_lines1") (fun () => { t_len = ##t })
    inl i', s'' = s |> advance_while ((=) '\n') t i
    if i' <> i
    then Ok (id, i', s'')
    else
        fun () =>
            inl preview_end = i + get_max_context () |> min s'.text_length
            "parsing.new_lines1 / expected at least one new line / "
            ++#? { rest = t |> slice i preview_end }
        |> Error
